module tb_top;

endmodule