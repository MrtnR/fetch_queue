package tb_package;

//`include "IFQ_if.sv"
`include "test1.sv"
`include "test2.sv"
`include "test3.sv"

endpackage