package tb_package;

//`include "IFQ_if.sv"
`include "test1.sv"

endpackage