module IFQ_ctrl(
    input clk,
    input reset,

    
)